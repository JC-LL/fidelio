fidelio_config_package_GCD.vhd